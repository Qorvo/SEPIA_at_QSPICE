* Zo_SEPIA0a.qsch
Rdcr N01 N03 2m
Cout DUTOUT N02 100�
Resr N02 0 2m
L1 N03 DUTOUT 50n
G1 0 DUTOUT CTRL 0 Istep
V2 CLK 0 PULSE 0 5 Tstep 1n 1n 0.5� 1�
شX1 �DUTOUT�d CLK�d� �CTRL�d o0�d o1�d� ��  SEPIA_v202 float Tstep={Tstep} float Tready={Tready} float Istep={Istep} char* Opt=vx
Iac 0 DUTOUT AC Iac
V1 N01 0 DC 5
* PyQSPICE TRAN begin
.param Iac = 0
.param Istep = -2
.param Tstep =  1mm
.param Tready = 0.9m 
.tran 2m
.plot tran V(dutout) V(o1)
.plot tran V(o0) 
* PyQSPICE TRAN end
* PyQSPICE AC begin
*.param Iac = 1
*.param Istep = 0
*.param Tstep =  999
*.param Tready = 998
*.ac dec 100 10 10Meg
*.plot ac V(out)
* PyQSPICE AC end
.end
